module tpu #()
()
endmodule